`include "light_rv32i_defs.vh"

module cpu_top (
    input wire clk,
    input wire reset   
);


    